module ABRO_blif(clk, rst, O, A, B, R);
input clk, rst;
output O;
input A;
input B;
input R;

wire A;
wire B;
wire R;
wire O;
wire w_0;
wire w_1;
wire R_O;
wire SM1_chk_0;
wire w_7;
wire w_8;
wire w_9;
wire SM3_chk_0;
wire w_10;
wire SM3_chk_1;
wire w_11;
wire SM10_chk_0;
wire w_12;
wire SM10_chk_1;
wire w_13;
wire B_O;
wire w_14;
wire w_15;
wire w_16;
wire w_17;
wire SM6_chk_0;
wire w_18;
wire SM6_chk_1;
wire w_19;
wire A_O;
wire w_20;
wire w_21;
wire w_22;
wire w_23;
wire w_24;
wire tick_O;
wire w_30;
wire w_31;
wire SM1_chk_1;
wire w_32;
wire SM1_goto_0;
wire SM1_goto_1;
wire SM1_hold;
wire w_36;
wire SM3_goto_0;
wire w_38;
wire SM3_goto_1;
wire SM3_hold;
wire SM6_goto_0;
wire w_42;
wire SM6_goto_1;
wire SM6_hold;
wire SM10_goto_0;
wire w_46;
wire SM10_goto_1;
wire SM10_hold;
wire ff_1_0_q;
wire ff_1_0_d;
wire g57;
wire ff_3_0_q;
wire ff_3_0_d;
wire g60;
wire ff_6_0_q;
wire ff_6_0_d;
wire g63;
wire ff_10_0_q;
wire ff_10_0_d;
wire g66;

assign O = w_24;
assign w_0 = 0;
assign w_1 = 1;
assign R_O = R;
assign SM1_chk_0 = !ff_1_0_q;
assign w_7 = R_O & SM1_chk_0;
assign w_8 = !R_O;
assign w_9 = w_8 & SM1_chk_0;
assign SM3_chk_0 = !ff_3_0_q;
assign w_10 = w_9 & SM3_chk_0;
assign SM3_chk_1 = ff_3_0_q;
assign w_11 = w_9 & SM3_chk_1;
assign SM10_chk_0 = !ff_10_0_q;
assign w_12 = w_11 & SM10_chk_0;
assign SM10_chk_1 = ff_10_0_q;
assign w_13 = w_11 & SM10_chk_1;
assign B_O = B;
assign w_14 = w_13 & B_O;
assign w_15 = !B_O;
assign w_16 = w_13 & w_15;
assign w_17 = w_14 | w_12;
assign SM6_chk_0 = !ff_6_0_q;
assign w_18 = w_11 & SM6_chk_0;
assign SM6_chk_1 = ff_6_0_q;
assign w_19 = w_11 & SM6_chk_1;
assign A_O = A;
assign w_20 = w_19 & A_O;
assign w_21 = !A_O;
assign w_22 = w_21 & w_19;
assign w_23 = w_20 | w_18;
assign w_24 = w_17 & w_23;
assign tick_O = w_1;
assign w_30 = !w_24;
assign w_31 = w_11 & w_30;
assign SM1_chk_1 = ff_1_0_q;
assign w_32 = w_9 | w_7 | SM1_chk_1;
assign SM1_goto_0 = w_32;
assign SM1_goto_1 = w_0;
assign SM1_hold = w_0;
assign w_36 = w_10 | w_24;
assign SM3_goto_0 = w_36;
assign w_38 = w_7 | w_31 | SM1_chk_1;
assign SM3_goto_1 = w_38;
assign SM3_hold = w_0;
assign SM6_goto_0 = w_23;
assign w_42 = w_7 | w_22 | SM1_chk_1;
assign SM6_goto_1 = w_42;
assign SM6_hold = w_0;
assign SM10_goto_0 = w_17;
assign w_46 = w_7 | w_16 | SM1_chk_1;
assign SM10_goto_1 = w_46;
assign SM10_hold = w_0;
d_ff1 u0(rst, clk, ff_1_0_q, ff_1_0_d);
assign ff_1_0_d = g57 | SM1_goto_1;
assign g57 = SM1_hold & ff_1_0_q;
d_ff0 u1(rst, clk, ff_3_0_q, ff_3_0_d);
assign ff_3_0_d = g60 | SM3_goto_1;
assign g60 = SM3_hold & ff_3_0_q;
d_ff0 u2(rst, clk, ff_6_0_q, ff_6_0_d);
assign ff_6_0_d = g63 | SM6_goto_1;
assign g63 = SM6_hold & ff_6_0_q;
d_ff0 u3(rst, clk, ff_10_0_q, ff_10_0_d);
assign ff_10_0_d = g66 | SM10_goto_1;
assign g66 = SM10_hold & ff_10_0_q;

endmodule
